library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use ieee.numeric_std.all;
use IEEE.STD_LOGIC_TEXTIO.ALL;
use std.textio.all;
entity Controller_tb is
end entity Controller_tb;

architecture behavioral of Controller_tb is

    -- Component Declaration for the memory
    component Memory
        Port ( Clk   : in  STD_LOGIC;
           Address : in  STD_LOGIC_VECTOR (7 downto 0);
           WriteEn : in  STD_LOGIC;
           DataIn  : in  STD_LOGIC_VECTOR (7 downto 0);
           DataOut    : out STD_LOGIC_VECTOR (7 downto 0));
    end component;

    -- Component Declaration for the Controller
    component Controller
        Port (
        Clk : in STD_LOGIC;
        Reset : in STD_LOGIC;
        Start,Lt : in STD_LOGIC;
        MaxWriteEn, MaxSrc, MinWriteEn, MinSrc, ValueWriteEn,IndexSrc, IndexWriteEn,AddrInWriteEn,AddrInSrc, AddressSrc, ALUOp : out STD_LOGIC;
        Done, ResultWriteEn : out STD_LOGIC;
        ALUSrcA, ALUSrcB : out std_logic_vector ( 1 downto 0)
    );
    end component;

    component Datapath
    PORT (Clk, Reset: IN STD_LOGIC;
          MaxWriteEn, MaxSrc, MinWriteEn, MinSrc, ValueWriteEn,
          IndexSrc, IndexWriteEn, AddrInWriteEn, AddrInSrc,
          AddressSrc, ALUOp: IN STD_LOGIC;
          ALUSrcA, ALUSrcB: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
          AddressIn, AddressOut, N, DataOut: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
          Lt: OUT STD_LOGIC;
          ALUResult, MemAddress: OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
	  TestMax,TestMin,TestValue,TestIdex,TestAddr: out STD_LOGIC_VECTOR (7 DOWNTO 0));
    end component;

    component Mux2
    GENERIC ( N : Integer := 8);
    Port (
        D0     : in  STD_LOGIC_VECTOR ( N - 1 downto 0);  -- Input A
        D1     : in  STD_LOGIC_VECTOR ( N - 1 downto 0);  -- Input B
        S   : in  STD_LOGIC;  -- Select signal
        Y     : out STD_LOGIC_VECTOR ( N - 1 downto 0)  -- Output Y
    );
    end component;

    component Mux1bit
    Port (
        D0     : in  STD_LOGIC;
        D1     : in  STD_LOGIC;
        S   : in  STD_LOGIC;  -- Select signal
        Y     : out STD_LOGIC
    );
    end component;

    -- Signals to connect to the memory component
    signal WriteEn     : std_logic := '0';
    signal Address   : std_logic_vector(7 downto 0) := (others => '0');
    signal DataIn  : std_logic_vector(7 downto 0) := (others => '0');
    signal DataOut : std_logic_vector(7 downto 0);
    file input_file : text open read_mode is "test.txt";
    file output_file : text open write_mode is "output.txt";

    signal Clk,Reset,Start,Lt    : std_logic := '0';
    signal MaxWriteEn, MaxSrc, MinWriteEn, MinSrc, ValueWriteEn,IndexSrc, IndexWriteEn,AddrInWriteEn,AddrInSrc, AddressSrc, ALUOp : std_logic:= '0';
    signal Done, ResultWriteEn : STD_LOGIC;
    signal ALUSrcA, ALUSrcB : std_logic_vector ( 1 downto 0);
    signal AddressIn,MemAddress,N,ALUResult,AddressOut : std_logic_vector(7 downto 0);
    signal TestMax,TestMin,TestValue,TestIdex,TestAddr: STD_LOGIC_VECTOR (7 DOWNTO 0);
    signal Select_Address_MemAddress: std_logic;
    signal output_mux: STD_LOGIC_VECTOR (7 DOWNTO 0);
    signal Select_Write_Enable: std_logic;
    signal output_mux2: std_logic;
    signal Select_DataIn : std_logic;
    signal output_datain_mux : std_logic_vector ( 7 downto 0);
    -- Function to convert std_logic_vector to string for display, dont need care about it
    function std_logic_vector_to_string(vector: std_logic_vector) return string is
        variable result : string(1 to vector'length);
    begin
        for i in vector'range loop
            if vector(i) = '1' then
                result(i+1) := '1';
            else
                result(i+1) := '0';
            end if;
        end loop;
        return result;
    end function;


    -- Clock period definition
    constant clk_period : time := 10 ns;
begin
   CTRL_UNIT: Controller
   Port map (
        Clk,
        Reset,
        Start,Lt,
        MaxWriteEn, MaxSrc, MinWriteEn, MinSrc, ValueWriteEn,IndexSrc, IndexWriteEn,AddrInWriteEn,AddrInSrc, AddressSrc, ALUOp,
        Done, ResultWriteEn,
        ALUSrcA,ALUSrcB
    );

   DATAPATH_UNIT: Datapath
   Port map (
	  Clk, Reset,
          MaxWriteEn, MaxSrc, MinWriteEn, MinSrc, ValueWriteEn,
          IndexSrc, IndexWriteEn, AddrInWriteEn, AddrInSrc,
          AddressSrc, ALUOp,
          ALUSrcA, ALUSrcB,
          AddressIn, AddressOut, N, DataOut,
          Lt,
          ALUResult, MemAddress,
	  TestMax,TestMin,TestValue,TestIdex,TestAddr
    );

    -- Instantiate the memory component
    MEMORY_UNIT: Memory
        port map (
            Clk    => Clk,
            WriteEn     => output_mux2,
            Address   => output_mux,
            DataIn  => output_datain_mux,
            DataOut => DataOut
        );

   address_Mux: Mux2
   Port map (
        Address,
	MemAddress,
	Select_Address_MemAddress,
	output_mux
    );

   Write_Enable_Mux: Mux1bit
   Port map (
        WriteEn,
	ResultWriteEn,
	Select_Write_Enable,
	output_mux2
    );

   DataIn_Mux: Mux2
   Port map (
        DataIn,
	ALUResult,
	Select_DataIn,
	output_datain_mux
    );
    -- Clock process definitions
    clk_process : process
    begin
        Clk <= '0';
        wait for clk_period/2;
        Clk <= '1';
        wait for clk_period/2;
    end process;

    -- Stimulus process
    stim_proc: process
	variable line_buffer : line;
	variable size: integer;
	variable data_buffer : std_logic_vector(7 downto 0);
	variable str : string(1 to 8);
    begin
	size:= 0;
	Select_DataIn <= '0';
	Select_Write_Enable <= '0';
	Select_Address_MemAddress <= '0';
	Address <= "00000000";
        -- Read lines from the file until end of file
        while not endfile(input_file) loop
            WriteEn <= '0';
            readline(input_file, line_buffer);
	    read(line_buffer, str);
             -- Convert string to std_logic_vector
            for i in 0 to 7 loop
                if str(i+1) = '0' then
                    data_buffer(7-i) := '0';
                elsif str(i+1) = '1' then
                    data_buffer(7-i) := '1';
                else
                    data_buffer(7-i) := '0'; -- Default case for non-binary characters
                end if;
            end loop;
	    report std_logic_vector_to_string(data_buffer);
	    size:= size + 1;
	    DataIn <= data_buffer;
	    WriteEn <= '1';
            wait until rising_edge(Clk);
	    Address <= Address + "00000001";
            -- Apply the data to the signal and wait for one clock cycle
        end loop;
        file_close(input_file);
	-- Compelete pushing all data from text file to memory
	
	Select_Address_MemAddress <= '1';
	WriteEn <= '0';
	AddressIn <= "00000000";
	AddressOut <= "01100100";
	--N <= "00001001";
	N <= std_logic_vector(to_unsigned(size, N'length));

	--Address <= MemAddress;
	wait for clk_period;
	wait for 2 ns;
        Start <= '1';
	--wait for 12*clk_period;
	--DataOut <= "10000000";
	wait until rising_edge(Done);
	Select_Write_Enable <= '1';
	Start <= '0';
	Select_DataIn <= '1'; 
	wait until rising_edge(Clk);
	Select_Write_Enable <= '0';
	WriteEn <= '0';
	wait for 2*clk_period;
	--Write to output.txt	
	write(line_buffer,std_logic_vector_to_string(DataOut));
	writeline(output_file,line_buffer);
	file_close(output_file);
	wait;
    end process;
end architecture behavioral;