LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_TEXTIO.ALL;
use std.textio.all;
ENTITY max_diff_tb IS
END ENTITY max_diff_tb;

ARCHITECTURE Behavioral OF max_diff_tb IS
    COMPONENT max_diff 
        Port ( Clk,Reset,Start   : in  STD_LOGIC;
               N,DataOut : in  STD_LOGIC_VECTOR (7 downto 0);
               AddressOut,AddressIn : in  STD_LOGIC_VECTOR (7 downto 0);
               Done ,ResultWriteEn: out  STD_LOGIC;
               MemAddress, ALUResult: out  STD_LOGIC_VECTOR (7 downto 0));
    END COMPONENT max_diff;
    COMPONENT Memory2 IS GENERIC (filename: STRING);
        PORT ( Clk   : IN  STD_LOGIC;
               Address : IN  STD_LOGIC_VECTOR (7 DOWNTO 0);
               WriteEn : IN  STD_LOGIC;
               DataIn  : IN  STD_LOGIC_VECTOR (7 DOWNTO 0);
               DataOut : OUT STD_LOGIC_VECTOR (7 DOWNTO 0));
    END COMPONENT Memory2;
    SIGNAL Clk, Reset, Start, Done, ResultWriteEn: STD_LOGIC;
    SIGNAL N, DataOut, AddressOut, AddressIn, MemAddress, ALUResult: STD_LOGIC_VECTOR (7 DOWNTO 0);
    CONSTANT clk_t: TIME := 10 NS;
    CONSTANT half_clk_t: TIME := clk_t / 2;
    file output_file : text open write_mode is "output.txt";

    -- Function to convert std_logic_vector to string for display, dont need care about it
    function std_logic_vector_to_string(vector: std_logic_vector) return string is
        variable result : string(1 to vector'length);
    begin
        for i in vector'range loop
            if vector(i) = '1' then
                result(9-(i+1)) := '1';
            else
                result(9-(i+1)) := '0';
            end if;
        end loop;
        return result;
    end function;

BEGIN
    dut: max_diff PORT MAP (Clk => Clk, Reset => Reset,
                    Start => Start, N => N, DataOut => DataOut,
                    AddressOut => AddressOut, AddressIn => AddressIn,
                    Done => Done, ResultWriteEn => ResultWriteEn,
                    MemAddress => MemAddress, ALUResult => ALUResult);
    memory_i: Memory2 GENERIC MAP (filename => "test.dat")
                      PORT MAP (Clk => Clk, Address => MemAddress,
                            WriteEn => ResultWriteEn, DataIn => ALUResult,
                            DataOut => DataOut);
                            
    PROCESS BEGIN
        Clk <= '0';
        WAIT FOR half_clk_t;
        Clk <= '1';
        WAIT FOR half_clk_t;
    END PROCESS;
    
    simu: PROCESS 
	variable line_buffer : line;
	BEGIN
        Reset <= '1';
        WAIT FOR clk_t;
        Reset <= '0';
        WAIT FOR clk_t / 10;
        Start <= '1';
        N <= "11111111";
        AddressIn <= "00000000";
        AddressOut <= "11111111";
        WAIT FOR 2 * clk_t;
        Start <= '0';
        
        WAIT UNTIL RISING_EDGE (Done);
	WAIT FOR clk_t;
	write(line_buffer,std_logic_vector_to_string(ALUResult));
        writeline(output_file,line_buffer);
   	file_close(output_file);
        WAIT;
    END PROCESS;
END ARCHITECTURE Behavioral;


